module int_ram#(
	parameter MEM_WIDTH = 8,
	parameter MEM_WORDS = 129
	) (
	input [$clog2(MEM_WORDS) - 1:0] address_1,
	input [$clog2(MEM_WORDS) - 1:0] address_2,
	input clk,
	input [MEM_WIDTH - 1:0] data_1,
	input [MEM_WIDTH - 1:0] data_2,
	input rden_1,
	input rden_2,
	input wren_1,
	input wren_2,
	output logic [MEM_WIDTH - 1:0] q_1,
	output logic [MEM_WIDTH - 1:0] q_2);

	altsyncram	altsyncram_component (
				.wren_a (wren_1),
				.clock0 (clk),
				.wren_b (wren_2),
				.address_a (address_1),
				.address_b (address_2),
				.rden_a (rden_1),
				.rden_b (rden_2),
				.data_a (data_1),
				.data_b (data_2),
				.q_a (q_1),
				.q_b (q_2),
				.aclr0 (1'b0),
				.aclr1 (1'b0),
				.addressstall_a (1'b0),
				.addressstall_b (1'b0),
				.byteena_a (1'b1),
				.byteena_b (1'b1),
				.clock1 (1'b1),
				.clocken0 (1'b1),
				.clocken1 (1'b1),
				.clocken2 (1'b1),
				.clocken3 (1'b1),
				.eccstatus ());
	defparam
		altsyncram_component.address_reg_b = "CLOCK0",
		altsyncram_component.clock_enable_input_a = "BYPASS",
		altsyncram_component.clock_enable_input_b = "BYPASS",
		altsyncram_component.clock_enable_output_a = "BYPASS",
		altsyncram_component.clock_enable_output_b = "BYPASS",
		altsyncram_component.indata_reg_b = "CLOCK0",
		altsyncram_component.intended_device_family = "Cyclone V",
		altsyncram_component.lpm_hint = "CLOCK_DUTY_CYCLE_DEPENDENCE=ON",
		altsyncram_component.lpm_type = "altsyncram",
		altsyncram_component.numwords_a = MEM_WORDS,
		altsyncram_component.numwords_b = MEM_WORDS,
		altsyncram_component.operation_mode = "BIDIR_DUAL_PORT",
		altsyncram_component.outdata_aclr_a = "NONE",
		altsyncram_component.outdata_aclr_b = "NONE",
		altsyncram_component.outdata_reg_a = "CLOCK0",
		altsyncram_component.outdata_reg_b = "CLOCK0",
		altsyncram_component.power_up_uninitialized = "FALSE",
		altsyncram_component.ram_block_type = "M10K",
		altsyncram_component.read_during_write_mode_mixed_ports = "OLD_DATA",
		altsyncram_component.read_during_write_mode_port_a = "NEW_DATA_NO_NBE_READ",
		altsyncram_component.read_during_write_mode_port_b = "NEW_DATA_NO_NBE_READ",
		altsyncram_component.widthad_a = $clog2(MEM_WORDS),
		altsyncram_component.widthad_b = $clog2(MEM_WORDS),
		altsyncram_component.width_a = MEM_WIDTH,
		altsyncram_component.width_b = MEM_WIDTH,
		altsyncram_component.width_byteena_a = 1,
		altsyncram_component.width_byteena_b = 1,
		altsyncram_component.wrcontrol_wraddress_reg_b = "CLOCK0";


endmodule